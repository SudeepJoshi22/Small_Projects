module mul2(
	input [2:0] a,
	output [3:0] y
);
assign y = a*2;

endmodule

module dff_const3(input clk, input reset, output reg q);
reg q1;

always @(posedge clk, posedge reset)
 begin
  if(reset) begin
   q <= 1'b1;
   q1 <= 1'b0;
  end
  else begin
   q1 <= 1'b1;
   q <= q1;
  end
 end
endmodule

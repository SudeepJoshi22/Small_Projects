module incomp_case (input i0 , input i1 , input i2 , input [1:0] sel, output reg y);
 always @ (*)
 begin
  case(sel)
   2'b00 : y = i0;
   2'b01 : y = i1;
  endcase
 end
endmodule

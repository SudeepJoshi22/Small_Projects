module dff_const2(input clk, input reset, output reg q);
 always @(posedge clk, posedge reset) begin
  if(reset)
   q <= 1'b1;
  else
   q <= 1'b1;
 end
endmodule

module incomp_if2 (input i0 , input i1 , input i2 , input i3, output reg y);
always @ (*)
 begin
  if(i0)
   y <= i1;
  else if (i2)
   y <= i3;

 end
endmodule

module partial_case_assign (input i0 , input i1 , input i2 , input [1:0] sel, output reg y , output reg x);
always @ (*)
begin
 case(sel)
  2'b00 : begin
   y = i0;
   x = i2;
   end
  2'b01 : y = i1;
  default : 
  begin
   x = i1;
   y = i2;
  end
 endcase
end
endmodule
